
module B;
import pkg::*;
initial
begin
#1;
no_of_trans=1;
#1;
display("From B");
end
endmodule
